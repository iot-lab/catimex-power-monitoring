* AD8539 SPICE Macro-model
* Description: Amplifier
* Generic Desc: 2.7/5V, CMOS, OP, Zero Drift, RRIO, 2X
* Developed by: ADISJ  HH
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (07/2010)
* Copyright 2007, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Node Assignments
*                  noninverting input
*                  |   inverting input
*                  |   |    positive supply
*                  |   |    |    negative supply
*                  |   |    |    |    output
*                  |   |    |    |    |
*                  |   |    |    |    |
.SUBCKT AD8539     1   2   99   50   45
*#ASSOC Category="Op-amps" symbol=opamp
*
* INPUT STAGE
*
M1  14  7  8  8 PIX L=1E-6 W=2.844E-05
M2  16  2  8  8 PIX L=1E-6 W=2.844E-05
M3  17  7 10 10 NIX L=1E-6 W=2.844E-05
M4  18  2 10 10 NIX L=1E-6 W=2.844E-05
RD1 14 50 2.667E+04
RD2 16 50 2.667E+04
RD3 99 17 2.667E+04
RD4 99 18 2.667E+04
C1  14 16 6.700E-12
C2  17 18 6.700E-12
I1  99  8 1.500E-05
I2  10 50 1.500E-05
V1  99  9 0.997E+00
V2  13 50 0.997E+00
D1   8  9 DX
D2  13 10 DX
EOS  7  1 POLY(4) (22,98) (73,98) (83,98) (70,98) 5.00E-06 1 1 1.2 1
IOS 1 2 1.00E-11
*
*CMRR=135dB, POLE AT 9 Hz ZERO AT 2.5 MHz
*
E1  21 98 POLY(2) (1,98) (2,98) 0 7.113E-02 7.113E-02
R10 21 22 1.592E+04
R20 22 98 1.989E-02
C10 21 22 1.000E-06
*
* PSRR=95dB, POLE AT 100 Hz
*
EPSY 72 98 POLY(1) (99,50) -8.89E-01 1.78E-00
CPS3 72 73 1.00E-06
RPS3 72 73 3.98E+04
RPS4 73 98 3.98E-02
*
* VOLTAGE NOISE REFERENCE OF 60nV/rt(Hz)
*
VN1 80 98 0
RN1 80 98  16.45E-05
*
HN  81 98 VN1 60E+00
RNHH1 81 183 5.3
CHH1 183 98 1uF
*
CHH2 183 184 2.7E-07
RNHH2 184 98 10
*
RNHH3 184 83 100k
CHH3 83 98 2.41E-10
*
* FLICKER NOISE CORNER = 0.000001 Hz
D5  69 98 DNOISE
VSN 69 98 DC 0.6551
H1  70 98 POLY(1) VSN 1.00E-03 1.00E+00
RN  70 98 1
*
* INTERNAL VOLTAGE REFERENCE
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) -242.5E-6 2.5E-06
EVP  97 98 POLY(1) (99,50) 0 0.5
EVN  51 98 POLY(1) (50,99) 0 0.5
*
* GAIN STAGE
G1 98 30 POLY(2) (14,16) (17,18) 0 2.678E-02 2.678E-02
R1 30 98 1.00E+06
V3 32 30 -3.603E-00
V4 30 33 -3.733E-00
EZ (145 0) (45 0) 1
CF 145 31 4.400E-08
RZ  30 31 3.800E+00
D3 32 97 DX
D4 51 33 DX
*
* OUTPUT STAGE
M5  45 46 99 99 POX L=1E-6 W=2.238E-05
M6  45 47 50 50 NOX L=1E-6 W=2.152E-05
EG1 99 46 POLY(1) (98,30) 1.299E+00 1
EG2 47 50 POLY(1) (30,98) 1.217E+00 1
*
* MODELS
.MODEL POX PMOS (LEVEL=2,KP=6.00E-05,VTO=-0.6,LAMBDA=0.02,RD=0)
.MODEL NOX NMOS (LEVEL=2,KP=8.00E-05,VTO=+0.6,LAMBDA=0.02,RD=0)
.MODEL PIX PMOS (LEVEL=2,KP=5.00E-05,VTO=-0.5,LAMBDA=0.02)
.MODEL NIX NMOS (LEVEL=2,KP=5.00E-05,VTO=0.5, LAMBDA=0.02)
.MODEL DX D(IS=1E-14,RS=5)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=2.50E-18)
*
.ENDS AD8539
*
*$




